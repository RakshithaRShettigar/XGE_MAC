`ifndef DESIGN_PKG_INCLUDED
`define DESIGN_PKG_INCLUDED

package design_pkg;





endpackage

`endif

