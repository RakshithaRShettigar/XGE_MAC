`ifndef DESIGN_PKG_OLD_INCLUDED_
`define DESIGN_PKG_OLD_INCLUDED_

package design_pkg_old;


`include "../rtl/fault_sm.sv"
`include "../rtl/generic_mem_small.sv"
`include "../rtl/generic_mem_medium.sv"
`include "../rtl/generic_fifo_ctrl.sv"
`include "../rtl/generic_fifo.sv"
`include "../rtl/meta_sync.sv"
`include "../rtl/meta_sync_single.sv"
`include "../rtl/rx_hold_fifo.sv"
`include "../rtl/rx_data_fifo.sv"
`include "../rtl/rx_dequeue.sv"
`include "../rtl/rx_enqueue.sv"
`include "../rtl/sync_clk_core.sv"
`include "../rtl/sync_clk_wb.sv"
`include "../rtl/sync_clk_xgmii_tx.sv"
`include "../rtl/tx_hold_fifo.sv"
`include "../rtl/tx_data_fifo.sv"
`include "../rtl/tx_dequeue.sv"
`include "../rtl/tx_enqueue.sv"
`include "../rtl/wishbone_if.sv"
`include "../rtl/xge_mac.sv"

  
endpackage

`endif
