shreyas
