`ifndef __XGEMAC_DEFINES_SV
`define __XGEMAC_DEFINES_SV

`define no_of_frames 8'd1

`endif
