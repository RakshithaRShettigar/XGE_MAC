ifndef AXI_ENV_PKG_INCLUDED_
`define AXI_ENV_PKG_INCLUDED_
package xgemac_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  //design

  

  


endpackage
